`timescale 1ns / 1ps
`include "aDefinitions.v"

////////////////////////////////////////////////////////////////////////////////////
//
// pGB, yet another FPGA fully functional and super fun GB classic clone!
// Copyright (C) 2015-2016  Diego Valverde (diego.valverde.g@gmail.com)
//
// This program is free software; you can redistribute it and/or
// modify it under the terms of the GNU General Public License
// as published by the Free Software Foundation; either version 2
// of the License, or (at your option) any later version.
//
// This program is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
//
// You should have received a copy of the GNU General Public License
// along with this program; if not, write to the Free Software
// Foundation, Inc., 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.
//
////////////////////////////////////////////////////////////////////////////////////
module pGB
(

input wire iClock,
input wire iReset

);

wire [15:0] wdZCPU_2_MMU_Addr;
wire [7:0]  wdZCPU_2_MMU_WriteData, wMMU_2_dzCPU_ReadData;
wire        wdZCPU_2_MMU_We;


mmu MMU
(
	.iClock( iClock ),
	.iReset( iReset ),
	.iCpuAddr(  wdZCPU_2_MMU_Addr ),
	.iWe(    wdZCPU_2_MMU_We   ),
	.iData(  wdZCPU_2_MMU_WriteData ),
	.oData(  wMMU_2_dzCPU_ReadData )
);

dzcpu  DZCPU
(
	.iClock( iClock ),
	.iReset( iReset ),
	.iMCUData( wMMU_2_dzCPU_ReadData ),
	.oMCUAddr( wdZCPU_2_MMU_Addr      ),
	.oMCUwe( wdZCPU_2_MMU_We ),
	.oMCUData( wdZCPU_2_MMU_WriteData )
);

endmodule
